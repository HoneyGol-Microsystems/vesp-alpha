module module_pwm #(

) (
    
);
    
endmodule