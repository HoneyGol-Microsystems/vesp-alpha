
module uart_top (
    input logic clk,
    input logic reset,
    input logic rx,

    output logic tx
);


endmodule