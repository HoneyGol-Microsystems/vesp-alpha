module pwm #(

) (
    
);
    
endmodule